// This is the unpowered netlist.
module user_proj_example (wb_clk_i,
    wb_rst_i,
    io_oeb,
    io_out);
 input wb_clk_i;
 input wb_rst_i;
 output [3:0] io_oeb;
 output [3:0] io_out;

 wire net6;
 wire net7;
 wire net8;
 wire net9;
 wire _00_;
 wire _01_;
 wire _02_;
 wire _03_;
 wire _04_;
 wire _05_;
 wire _06_;
 wire _07_;
 wire _08_;
 wire clknet_0_wb_clk_i;
 wire clknet_1_0__leaf_wb_clk_i;
 wire clknet_1_1__leaf_wb_clk_i;
 wire net1;
 wire net10;
 wire net11;
 wire net12;
 wire net13;
 wire net14;
 wire net15;
 wire net16;
 wire net17;
 wire net2;
 wire net3;
 wire net4;
 wire net5;

 sky130_fd_sc_hd__diode_2 ANTENNA_hold2_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_hold6_A (.DIODE(net5));
 sky130_fd_sc_hd__diode_2 ANTENNA_output4_A (.DIODE(net4));
 sky130_fd_sc_hd__diode_2 ANTENNA_output5_A (.DIODE(net5));
 sky130_fd_sc_hd__decap_3 FILLER_0_0_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_0_141 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_154 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_0_166 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_0_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_0_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_0_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_10_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_157 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_10_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_10_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_10_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_137 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_11_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_11_157 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_163 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_11_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_187 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_11_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_11_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_11_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_12_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_12_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_12_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_13_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_13_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_13_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_13_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_14_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_14_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_14_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_15_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_15_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_15_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_15_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_15_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_16_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_16_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_16_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_17_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_17_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_17_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_17_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_17_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_18_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_18_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_18_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_19_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_19_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_19_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_19_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_19_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_1_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_161 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_1_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_1_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_1_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_20_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_20_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_20_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_21_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_21_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_21_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_21_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_21_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_22_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_22_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_22_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_23_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_23_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_23_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_23_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_23_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_24_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_24_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_24_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_25_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_25_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_25_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_25_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_26_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_26_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_26_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_27_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_27_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_27_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_27_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_27_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_28_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_28_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_28_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_29_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_29_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_29_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_29_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_29_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_2_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_157 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_2_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_2_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_2_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_30_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_30_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_30_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_31_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_31_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_31_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_31_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_31_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_32_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_32_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_32_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_33_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_33_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_33_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_33_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_33_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_34_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_34_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_34_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_35_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_35_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_35_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_35_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_35_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_36_177 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_36_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_36_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_36_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_36_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_37_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_37_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_37_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_37_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_37_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_38_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_38_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_38_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_39_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_39_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_39_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_39_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_39_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_3_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_15 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_3_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_3_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_3_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_40_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_40_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_40_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_41_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_41_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_41_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_41_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_41_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_42_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_42_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_42_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_43_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_43_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_43_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_43_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_43_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_44_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_44_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_44_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_45_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_45_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_45_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_45_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_45_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_46_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_46_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_46_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_47_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_47_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_47_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_47_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_47_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_153 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_171 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_48_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_48_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_48_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_49_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_49_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_49_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_49_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_49_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_153 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_4_186 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_4_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_4_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_4_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_50_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_50_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_50_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_51_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_51_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_51_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_51_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_51_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_52_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_52_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_52_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_53_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_53_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_53_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_53_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_53_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_54_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_54_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_54_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_55_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_55_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_55_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_55_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_55_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_56_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_56_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_56_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_57_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_57_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_57_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_57_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_57_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_58_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_58_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_58_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_59_181 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_59_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_59_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_59_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_5_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_15 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_5_165 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_5_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_5_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_5_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_60_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_60_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_60_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_61_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_61_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_61_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_61_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_61_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_62_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_62_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_62_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_63_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_63_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_63_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_63_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_63_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_64_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_64_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_64_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_65_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_65_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_65_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_65_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_65_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_66_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_66_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_66_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_67_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_67_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_67_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_67_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_67_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_68_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_68_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_68_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_69_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_69_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_69_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_69_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_69_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_15 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_6_153 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_157 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_178 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_6_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_6_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_6_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_165 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_70_177 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_70_185 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_70_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_70_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_70_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_71_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_167 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_173 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_71_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_71_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_71_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_72_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_72_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_72_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_73_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_73_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_73_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_73_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_73_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_74_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_74_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_74_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_75_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_75_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_75_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_75_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_75_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_76_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_76_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_76_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_77_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_77_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_77_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_77_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_77_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_78_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_78_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_78_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_79_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_79_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_79_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_79_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_79_93 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_7_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_7_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_7_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_7_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_7_93 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_153 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_177 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_189 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_80_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_80_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_80_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_15 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_81_161 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_167 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_169 ();
 sky130_fd_sc_hd__decap_8 FILLER_0_81_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_81_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_81_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_81_93 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_125 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_137 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_15 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_165 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_169 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_82_181 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_82_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_41 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_69 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_82_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_82_97 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_109 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_121 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_133 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_139 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_141 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_8_153 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_8_187 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_29 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_41 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_53 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_65 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_8_77 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_8_83 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_85 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_8_97 ();
 sky130_fd_sc_hd__decap_6 FILLER_0_9_105 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_111 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_113 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_125 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_137 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_149 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_15 ();
 sky130_fd_sc_hd__fill_2 FILLER_0_9_166 ();
 sky130_fd_sc_hd__decap_3 FILLER_0_9_169 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_189 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_27 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_3 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_39 ();
 sky130_fd_sc_hd__decap_4 FILLER_0_9_51 ();
 sky130_fd_sc_hd__fill_1 FILLER_0_9_55 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_57 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_69 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_81 ();
 sky130_ef_sc_hd__decap_12 FILLER_0_9_93 ();
 sky130_fd_sc_hd__decap_3 PHY_0 ();
 sky130_fd_sc_hd__decap_3 PHY_1 ();
 sky130_fd_sc_hd__decap_3 PHY_10 ();
 sky130_fd_sc_hd__decap_3 PHY_100 ();
 sky130_fd_sc_hd__decap_3 PHY_101 ();
 sky130_fd_sc_hd__decap_3 PHY_102 ();
 sky130_fd_sc_hd__decap_3 PHY_103 ();
 sky130_fd_sc_hd__decap_3 PHY_104 ();
 sky130_fd_sc_hd__decap_3 PHY_105 ();
 sky130_fd_sc_hd__decap_3 PHY_106 ();
 sky130_fd_sc_hd__decap_3 PHY_107 ();
 sky130_fd_sc_hd__decap_3 PHY_108 ();
 sky130_fd_sc_hd__decap_3 PHY_109 ();
 sky130_fd_sc_hd__decap_3 PHY_11 ();
 sky130_fd_sc_hd__decap_3 PHY_110 ();
 sky130_fd_sc_hd__decap_3 PHY_111 ();
 sky130_fd_sc_hd__decap_3 PHY_112 ();
 sky130_fd_sc_hd__decap_3 PHY_113 ();
 sky130_fd_sc_hd__decap_3 PHY_114 ();
 sky130_fd_sc_hd__decap_3 PHY_115 ();
 sky130_fd_sc_hd__decap_3 PHY_116 ();
 sky130_fd_sc_hd__decap_3 PHY_117 ();
 sky130_fd_sc_hd__decap_3 PHY_118 ();
 sky130_fd_sc_hd__decap_3 PHY_119 ();
 sky130_fd_sc_hd__decap_3 PHY_12 ();
 sky130_fd_sc_hd__decap_3 PHY_120 ();
 sky130_fd_sc_hd__decap_3 PHY_121 ();
 sky130_fd_sc_hd__decap_3 PHY_122 ();
 sky130_fd_sc_hd__decap_3 PHY_123 ();
 sky130_fd_sc_hd__decap_3 PHY_124 ();
 sky130_fd_sc_hd__decap_3 PHY_125 ();
 sky130_fd_sc_hd__decap_3 PHY_126 ();
 sky130_fd_sc_hd__decap_3 PHY_127 ();
 sky130_fd_sc_hd__decap_3 PHY_128 ();
 sky130_fd_sc_hd__decap_3 PHY_129 ();
 sky130_fd_sc_hd__decap_3 PHY_13 ();
 sky130_fd_sc_hd__decap_3 PHY_130 ();
 sky130_fd_sc_hd__decap_3 PHY_131 ();
 sky130_fd_sc_hd__decap_3 PHY_132 ();
 sky130_fd_sc_hd__decap_3 PHY_133 ();
 sky130_fd_sc_hd__decap_3 PHY_134 ();
 sky130_fd_sc_hd__decap_3 PHY_135 ();
 sky130_fd_sc_hd__decap_3 PHY_136 ();
 sky130_fd_sc_hd__decap_3 PHY_137 ();
 sky130_fd_sc_hd__decap_3 PHY_138 ();
 sky130_fd_sc_hd__decap_3 PHY_139 ();
 sky130_fd_sc_hd__decap_3 PHY_14 ();
 sky130_fd_sc_hd__decap_3 PHY_140 ();
 sky130_fd_sc_hd__decap_3 PHY_141 ();
 sky130_fd_sc_hd__decap_3 PHY_142 ();
 sky130_fd_sc_hd__decap_3 PHY_143 ();
 sky130_fd_sc_hd__decap_3 PHY_144 ();
 sky130_fd_sc_hd__decap_3 PHY_145 ();
 sky130_fd_sc_hd__decap_3 PHY_146 ();
 sky130_fd_sc_hd__decap_3 PHY_147 ();
 sky130_fd_sc_hd__decap_3 PHY_148 ();
 sky130_fd_sc_hd__decap_3 PHY_149 ();
 sky130_fd_sc_hd__decap_3 PHY_15 ();
 sky130_fd_sc_hd__decap_3 PHY_150 ();
 sky130_fd_sc_hd__decap_3 PHY_151 ();
 sky130_fd_sc_hd__decap_3 PHY_152 ();
 sky130_fd_sc_hd__decap_3 PHY_153 ();
 sky130_fd_sc_hd__decap_3 PHY_154 ();
 sky130_fd_sc_hd__decap_3 PHY_155 ();
 sky130_fd_sc_hd__decap_3 PHY_156 ();
 sky130_fd_sc_hd__decap_3 PHY_157 ();
 sky130_fd_sc_hd__decap_3 PHY_158 ();
 sky130_fd_sc_hd__decap_3 PHY_159 ();
 sky130_fd_sc_hd__decap_3 PHY_16 ();
 sky130_fd_sc_hd__decap_3 PHY_160 ();
 sky130_fd_sc_hd__decap_3 PHY_161 ();
 sky130_fd_sc_hd__decap_3 PHY_162 ();
 sky130_fd_sc_hd__decap_3 PHY_163 ();
 sky130_fd_sc_hd__decap_3 PHY_164 ();
 sky130_fd_sc_hd__decap_3 PHY_165 ();
 sky130_fd_sc_hd__decap_3 PHY_17 ();
 sky130_fd_sc_hd__decap_3 PHY_18 ();
 sky130_fd_sc_hd__decap_3 PHY_19 ();
 sky130_fd_sc_hd__decap_3 PHY_2 ();
 sky130_fd_sc_hd__decap_3 PHY_20 ();
 sky130_fd_sc_hd__decap_3 PHY_21 ();
 sky130_fd_sc_hd__decap_3 PHY_22 ();
 sky130_fd_sc_hd__decap_3 PHY_23 ();
 sky130_fd_sc_hd__decap_3 PHY_24 ();
 sky130_fd_sc_hd__decap_3 PHY_25 ();
 sky130_fd_sc_hd__decap_3 PHY_26 ();
 sky130_fd_sc_hd__decap_3 PHY_27 ();
 sky130_fd_sc_hd__decap_3 PHY_28 ();
 sky130_fd_sc_hd__decap_3 PHY_29 ();
 sky130_fd_sc_hd__decap_3 PHY_3 ();
 sky130_fd_sc_hd__decap_3 PHY_30 ();
 sky130_fd_sc_hd__decap_3 PHY_31 ();
 sky130_fd_sc_hd__decap_3 PHY_32 ();
 sky130_fd_sc_hd__decap_3 PHY_33 ();
 sky130_fd_sc_hd__decap_3 PHY_34 ();
 sky130_fd_sc_hd__decap_3 PHY_35 ();
 sky130_fd_sc_hd__decap_3 PHY_36 ();
 sky130_fd_sc_hd__decap_3 PHY_37 ();
 sky130_fd_sc_hd__decap_3 PHY_38 ();
 sky130_fd_sc_hd__decap_3 PHY_39 ();
 sky130_fd_sc_hd__decap_3 PHY_4 ();
 sky130_fd_sc_hd__decap_3 PHY_40 ();
 sky130_fd_sc_hd__decap_3 PHY_41 ();
 sky130_fd_sc_hd__decap_3 PHY_42 ();
 sky130_fd_sc_hd__decap_3 PHY_43 ();
 sky130_fd_sc_hd__decap_3 PHY_44 ();
 sky130_fd_sc_hd__decap_3 PHY_45 ();
 sky130_fd_sc_hd__decap_3 PHY_46 ();
 sky130_fd_sc_hd__decap_3 PHY_47 ();
 sky130_fd_sc_hd__decap_3 PHY_48 ();
 sky130_fd_sc_hd__decap_3 PHY_49 ();
 sky130_fd_sc_hd__decap_3 PHY_5 ();
 sky130_fd_sc_hd__decap_3 PHY_50 ();
 sky130_fd_sc_hd__decap_3 PHY_51 ();
 sky130_fd_sc_hd__decap_3 PHY_52 ();
 sky130_fd_sc_hd__decap_3 PHY_53 ();
 sky130_fd_sc_hd__decap_3 PHY_54 ();
 sky130_fd_sc_hd__decap_3 PHY_55 ();
 sky130_fd_sc_hd__decap_3 PHY_56 ();
 sky130_fd_sc_hd__decap_3 PHY_57 ();
 sky130_fd_sc_hd__decap_3 PHY_58 ();
 sky130_fd_sc_hd__decap_3 PHY_59 ();
 sky130_fd_sc_hd__decap_3 PHY_6 ();
 sky130_fd_sc_hd__decap_3 PHY_60 ();
 sky130_fd_sc_hd__decap_3 PHY_61 ();
 sky130_fd_sc_hd__decap_3 PHY_62 ();
 sky130_fd_sc_hd__decap_3 PHY_63 ();
 sky130_fd_sc_hd__decap_3 PHY_64 ();
 sky130_fd_sc_hd__decap_3 PHY_65 ();
 sky130_fd_sc_hd__decap_3 PHY_66 ();
 sky130_fd_sc_hd__decap_3 PHY_67 ();
 sky130_fd_sc_hd__decap_3 PHY_68 ();
 sky130_fd_sc_hd__decap_3 PHY_69 ();
 sky130_fd_sc_hd__decap_3 PHY_7 ();
 sky130_fd_sc_hd__decap_3 PHY_70 ();
 sky130_fd_sc_hd__decap_3 PHY_71 ();
 sky130_fd_sc_hd__decap_3 PHY_72 ();
 sky130_fd_sc_hd__decap_3 PHY_73 ();
 sky130_fd_sc_hd__decap_3 PHY_74 ();
 sky130_fd_sc_hd__decap_3 PHY_75 ();
 sky130_fd_sc_hd__decap_3 PHY_76 ();
 sky130_fd_sc_hd__decap_3 PHY_77 ();
 sky130_fd_sc_hd__decap_3 PHY_78 ();
 sky130_fd_sc_hd__decap_3 PHY_79 ();
 sky130_fd_sc_hd__decap_3 PHY_8 ();
 sky130_fd_sc_hd__decap_3 PHY_80 ();
 sky130_fd_sc_hd__decap_3 PHY_81 ();
 sky130_fd_sc_hd__decap_3 PHY_82 ();
 sky130_fd_sc_hd__decap_3 PHY_83 ();
 sky130_fd_sc_hd__decap_3 PHY_84 ();
 sky130_fd_sc_hd__decap_3 PHY_85 ();
 sky130_fd_sc_hd__decap_3 PHY_86 ();
 sky130_fd_sc_hd__decap_3 PHY_87 ();
 sky130_fd_sc_hd__decap_3 PHY_88 ();
 sky130_fd_sc_hd__decap_3 PHY_89 ();
 sky130_fd_sc_hd__decap_3 PHY_9 ();
 sky130_fd_sc_hd__decap_3 PHY_90 ();
 sky130_fd_sc_hd__decap_3 PHY_91 ();
 sky130_fd_sc_hd__decap_3 PHY_92 ();
 sky130_fd_sc_hd__decap_3 PHY_93 ();
 sky130_fd_sc_hd__decap_3 PHY_94 ();
 sky130_fd_sc_hd__decap_3 PHY_95 ();
 sky130_fd_sc_hd__decap_3 PHY_96 ();
 sky130_fd_sc_hd__decap_3 PHY_97 ();
 sky130_fd_sc_hd__decap_3 PHY_98 ();
 sky130_fd_sc_hd__decap_3 PHY_99 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_166 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_167 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_168 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_169 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_170 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_171 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_172 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_173 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_174 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_175 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_176 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_177 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_178 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_179 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_180 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_181 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_182 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_183 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_184 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_185 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_186 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_187 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_188 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_189 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_190 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_191 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_192 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_193 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_194 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_195 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_196 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_197 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_198 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_199 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_200 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_201 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_202 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_203 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_204 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_205 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_206 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_207 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_208 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_209 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_210 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_211 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_212 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_213 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_214 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_215 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_216 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_217 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_218 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_219 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_220 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_221 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_222 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_223 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_224 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_225 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_226 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_227 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_228 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_229 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_230 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_231 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_232 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_233 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_234 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_235 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_236 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_237 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_238 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_239 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_240 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_241 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_242 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_243 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_244 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_245 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_246 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_247 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_248 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_249 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_250 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_251 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_252 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_253 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_254 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_255 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_256 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_257 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_258 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_259 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_260 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_261 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_262 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_263 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_264 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_265 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_266 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_267 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_268 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_269 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_270 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_271 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_272 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_273 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_274 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_275 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_276 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_277 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_278 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_279 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_280 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_281 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_282 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_283 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_284 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_285 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_286 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_287 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_288 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_289 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_290 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_291 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_292 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_293 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_294 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_295 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_296 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_297 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_298 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_299 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_300 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_301 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_302 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_303 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_304 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_305 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_306 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_307 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_308 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_309 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_310 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_311 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_312 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_313 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_314 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_315 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_316 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_317 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_318 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_319 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_320 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_321 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_322 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_323 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_324 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_325 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_326 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_327 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_328 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_329 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_330 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_331 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_332 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_333 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_334 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_335 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_336 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_337 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_338 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_339 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_340 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_341 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_342 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_343 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_344 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_345 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_346 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_347 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_348 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_349 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_350 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_351 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_352 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_353 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_354 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_355 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_356 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_357 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_358 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_359 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_360 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_361 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_362 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_363 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_364 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_365 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_366 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_367 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_368 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_369 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_370 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_371 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_372 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_373 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_374 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_375 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_376 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_377 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_378 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_379 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_380 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_381 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_382 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_383 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_384 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_385 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_386 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_387 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_388 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_389 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_390 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_391 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_392 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_393 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_394 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_395 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_396 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_397 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_398 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_399 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_400 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_401 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_402 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_403 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_404 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_405 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_406 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_407 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_408 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_409 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_410 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_411 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_412 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_413 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_414 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_415 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_416 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_417 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_418 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_419 ();
 sky130_fd_sc_hd__tapvpwrvgnd_1 TAP_420 ();
 sky130_fd_sc_hd__nor2_1 _09_ (.A(net10),
    .B(net1),
    .Y(_00_));
 sky130_fd_sc_hd__a21oi_1 _10_ (.A1(net10),
    .A2(net14),
    .B1(net1),
    .Y(_04_));
 sky130_fd_sc_hd__o21a_1 _11_ (.A1(net10),
    .A2(net14),
    .B1(_04_),
    .X(_01_));
 sky130_fd_sc_hd__a21oi_1 _12_ (.A1(net10),
    .A2(net3),
    .B1(net11),
    .Y(_05_));
 sky130_fd_sc_hd__a31o_1 _13_ (.A1(net10),
    .A2(net3),
    .A3(net11),
    .B1(net1),
    .X(_06_));
 sky130_fd_sc_hd__nor2_1 _14_ (.A(net12),
    .B(_06_),
    .Y(_02_));
 sky130_fd_sc_hd__nand4_1 _15_ (.A(net10),
    .B(net14),
    .C(net11),
    .D(net15),
    .Y(_07_));
 sky130_fd_sc_hd__a31o_1 _16_ (.A1(net10),
    .A2(net14),
    .A3(net11),
    .B1(net15),
    .X(_08_));
 sky130_fd_sc_hd__and3b_1 _17_ (.A_N(net1),
    .B(_07_),
    .C(_08_),
    .X(_03_));
 sky130_fd_sc_hd__dfxtp_1 _18_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_00_),
    .Q(net2));
 sky130_fd_sc_hd__dfxtp_2 _19_ (.CLK(clknet_1_0__leaf_wb_clk_i),
    .D(_01_),
    .Q(net3));
 sky130_fd_sc_hd__dfxtp_1 _20_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(net13),
    .Q(net4));
 sky130_fd_sc_hd__dfxtp_2 _21_ (.CLK(clknet_1_1__leaf_wb_clk_i),
    .D(_03_),
    .Q(net5));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_0_wb_clk_i (.A(wb_clk_i),
    .X(clknet_0_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_0__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_0__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_16 clkbuf_1_1__f_wb_clk_i (.A(clknet_0_wb_clk_i),
    .X(clknet_1_1__leaf_wb_clk_i));
 sky130_fd_sc_hd__clkbuf_2 hold1 (.A(net16),
    .X(net10));
 sky130_fd_sc_hd__buf_1 hold2 (.A(net4),
    .X(net11));
 sky130_fd_sc_hd__dlygate4sd3_1 hold3 (.A(_05_),
    .X(net12));
 sky130_fd_sc_hd__dlygate4sd3_1 hold4 (.A(_02_),
    .X(net13));
 sky130_fd_sc_hd__dlymetal6s2s_1 hold5 (.A(net17),
    .X(net14));
 sky130_fd_sc_hd__dlygate4sd3_1 hold6 (.A(net5),
    .X(net15));
 sky130_fd_sc_hd__dlygate4sd3_1 hold7 (.A(net2),
    .X(net16));
 sky130_fd_sc_hd__dlygate4sd3_1 hold8 (.A(net3),
    .X(net17));
 sky130_fd_sc_hd__buf_1 input1 (.A(wb_rst_i),
    .X(net1));
 sky130_fd_sc_hd__buf_12 output2 (.A(net2),
    .X(io_out[0]));
 sky130_fd_sc_hd__buf_12 output3 (.A(net3),
    .X(io_out[1]));
 sky130_fd_sc_hd__buf_12 output4 (.A(net4),
    .X(io_out[2]));
 sky130_fd_sc_hd__buf_12 output5 (.A(net5),
    .X(io_out[3]));
 sky130_fd_sc_hd__conb_1 user_proj_example_6 (.LO(net6));
 sky130_fd_sc_hd__conb_1 user_proj_example_7 (.LO(net7));
 sky130_fd_sc_hd__conb_1 user_proj_example_8 (.LO(net8));
 sky130_fd_sc_hd__conb_1 user_proj_example_9 (.LO(net9));
 assign io_oeb[0] = net6;
 assign io_oeb[1] = net7;
 assign io_oeb[2] = net8;
 assign io_oeb[3] = net9;
endmodule

